module sr_ff(
    input  wire clk,
    input  wire s,
    input  wire r,
    output reg  q,
    output wire nq
);
    always @(posedge clk) begin
        case ({s, r})
            2'b10: q <= 1'b1;
            2'b01: q <= 1'b0;
            2'b00: q <= q;
            2'b11: q <= 1'bx;
        endcase
    end
    assign nq = ~q;
endmodule